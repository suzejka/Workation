��        �sklearn.linear_model._ridge��Ridge���)��}�(�alpha�G?�      �fit_intercept���	normalize���copy_X���max_iter�N�tol�G?PbM����solver��auto��random_state�M��n_features_in_�M��coef_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KM���h�dtype����f4�����R�(K�<�NNNJ����J����K t�b�B�   ;���6���D��D���}���bEK������/n��yf�ľR�C83���e�"K�E]_#ƅR?�2�FVO;���D�D4��E�K1ŮG_��,E    �d�a��D]���@�D���mEjGE��E�cE�����1���F    (i���rE>5OŎ�mĔ�ŒeDشVE����B��E���x�Ƶ�;�.ZJE    HCA�$*EE�E'E�ϰ�    �eV�u�ES�D�ͨ��Zť��[��Z��Ej^�Dn��Ea
 E���D�#�-���{�D�T�ŗS�D)(�E��7D?�+ElߥD�+�E�X�E�Q+�gE���E3'DF˓ů�bEa����RT�u�!ďX�E�B��k��� F�N����Exrwž���f����7EW�� %�M9pE���D��'E�~�Ŵ�Dt�tE�n#�'F$E�DyE6������+�uE/;����F� �D�q��L҄ś�Ďs�ě!GEɒ�=��&1�ň�EZ�[�8L�D��:Ci0�E]��C3 Cź�&�_��DQ�#��0�{'fE;�}�    �.�D��Ũ�E���Ŗx�DL@����EԶQ�+=2EHq7E��E��DZ���ZH��y�d��.Cv�H�*%��!ԗE��E        ���y�c�#D    �+�D�֭D�
œlSE�R|ę������        ���Ŀ��DI�����%����-E (D���C    ���B8-��EK�D��8�0�E    )6�y���F)�
E������z���葮D    A��D�#�        ƊFE    ̡�Ī��(�    vy�            j>��@Կ�    8a"Ð�Kł��DR�`E�ע�3��            |]�Ci��D��C^ܢ�5-E    ��Er/x�    ��#ůw7E���C���D        �~�����    A�2E�"�Ė6�E    �J�    K �E    �0mEl�D�q��        ��kE�/�E�I�ık�Do�pE    ��eŷp�D��!E�A�D���E��LE��E<�Djf�Ķ�E5�D	:C�ҋ�H�	�-!cE��XE��lF-/;D��E>�%�|�'�{�D��p����    �S�E�R�Ā�D��<��+�H�0�f�C��}�    �H�Eq9[E�D ��ݶsE    =s#�ű�EEs�E    ���    ���D���E���C�E�[j�&�DO	��)5�DwgE    [�GE��jĿaEd|oœN4�    
;ŵQE9g]E�'?E�>���>Dk���:�D    *��D�uxD����    �*���|(E    ���Dav���JD�    /75E�p��V�V�    ۣ�Ĩ�(� 9Eʂ�C    �K�Ĩ��DZ%��ol�D ���            ���şgO�0�;�b��;�\]�    �R�D唝�                ��IE�����ZE*�E    ��s�8��XP�C�2�� RE        w�CɃ��?��    �f�O�
D��cŲ��D*�8D.�lE3���*ސD��h�FҵC    kc*�q����!zD"F@^JE+��ÿ��x��!FE���:#�Â��DHl�D���;gxă�G��Ek'�E|щC��D»��v�ĕ	:Ţl[�    hDR�C�    �D"��PģX���E܍E�l�A3��jP��;:[���E    x0��N(E    ���Bj��K�        1�+,E�K�ܠ�D��D���B�.2C            I��DP��D�H��    ۭ�ĕ�5�G���!�    �	��@��ك_E>���        u|�EDt�D�o���?�D	��C�uD    �%C    L�Ej gD��gğA�D��Dč�D�=s	E�?��!���}4E��DZ�Ch�|DO%D��CEn�cE�:�C�^��krCE    �ǾD���o���f�E��Āp�D�U�Ä��ĝAfE    ۄJŶ,WE�=�ä�Ū}PD        ���        ��JţCjM�DUY�f����OP�c��B        u����E    �<D�����DE            ����    �L����    �k~D����    &��37�D    �pŗ [�83�C��?�        �22Dm�D��    �$���FE�`�        �{��݄Ğ2��V#�Cµ&C        �|D�[CC�8�uA�E���D�C�Ej�kE    37�D��&Ş;5E�X��        ���"��D��ᒞE���ė��İ�D    3�<E������T�Zֻ�
#D�~'DLԄD�E���D�9E    ��0�        u���    6��D        ��D][-F�zFdi�D$j�C        O`�E��;E    a���rT�D��B����_��\ec�Q�OE�^��B�Ă�EQ4�DP���E����    ��E���A    =[đ�Z�A��DG�����F�_%C    rL��    V�lĩ���;���ElŎ�+�    (�D��B�������+���e�     �E    Z�DvnE����Hq�E    >��C�*�h�2űd+Dnm�D    �� Eq��E�Y��        +Q#�sD    �fD�
E�͊D��"EE}�)�        �(E��eEu ��`WD�ҽD	���cEL'E�6�D~��-�D�GF+�$EE�DSqpC/��    ��C    ���D�b�D�˵D�3��ύ�E!Q{E�y�D*;��8�=F%#�D    VH�ú��    Dd�Ń���W��CQ�i�    ��sE��Ŷ��C�E[�E    �k�E��ID��F�%SŨ� �    �H$EﳛEz�.�\�E����%�&C�I%�    <�g�e�v�!�Dp0�ĻE����VX��bŕs�F��'F    ���E���DՇ�C6VEt�8E�8�E    �"P��7E���A    ��E$�ĺA�ŴC]�����w�o�O�~Q�D�~�Đ�kĶ �C�t�E    6�rĩ{@��7g���D��D�į7��    '��D=��C݅��s�D�����*�D�-��>^�gt�        ��l� ��D���        G2��M��~v�����,}D�(�C	��+kEWE            �
�    �x1E�����;D9��D    �1ű�JE    �w�E�)JķV�(��F�82ƕdų��EJ&EQѰ�)���P�E        ��ź_D(-fE�ky�rN�7�EwvPE���E�F�N�D�v���a�Em D    c��ݬ�    � C�_�ðs�E��|�    s�ELiG�    �<E�ȶD�ǵD    -/�F�LE\HE    ��>D�dF    ʖ&F�@MF��Efp�C����S-EXHh�zK8�ZX�-�m�(à���DgA�{��DRC@���G��C    ��	E���E_@YF    �	�;�Ct�D F��8��E�>9E��E    �@EI�_�`P=D    �3E��E�4e��    Q�D���ßǓD�.}C� ?����    �PL�C�ƇD%{�Eg�|E]z9� �iĴZ�C    �C��    ��DO@E��_Ez��1f}E��$E    YD��ND    �z�D���z}��hE8�ā��D�ҴD��t�H�7E    ��A���        �E�            &:"E��nD�����d���h�D���C��P�*)�}YqE                :�E�( E�V�D�!��81ń���H`-E���D��Dt���+^E    �4����TDBkw�,���Җ��cA��>]�Ö-E            s����f��    ���D[Z�D{�s�n�
��4E    }%�F�?Ń�|F�        �{8�Ȥ!D    ��ķw&����n�D    H��E)ٚDu�0���Xň�D�f��ͻ�        ���8y1����DQ&�E�ߵD�۳D�&�    ��F�e��    ���    ��Fv��F�^?�    2p�Mw�Eg�D    ���C    �H4F    7�&F�"F��)�P=#F���E,�ZF    ӕ��    $�F
0��    �$F���0�qB����gYFy��E �Dq��    �+v�    )�dF�~S��@��`EK�M��9ů�Dd�E�DXD_��s�>���D�+DC<�Cq_�DJ������8����3C�'w�c>�B� �7
pE�-�D�ҺC
�Y�v�/Dm��D�ϘDԤ4EV�� �/D��>����2Eb���E��R�D���E��T%ZĞ@KC�P�ƫCE:D��^��DS6�D����@��uEL������qyãW�D�QTŉǒEk]Ĥb�$��C�ŚD+��Dϡ�Df�@ĝ��EyQ�@S��%�C�S��t �a
Ep���� ��D���n�.D                �BC���"D� O�~{������?��C�L7�a�M�V9�    ,���|�D    !�    ��ŧȮ�Sa���j=D��}D    ����        ��Ľ���g��p?D���D{ :ā�%E�C�������D��ʹ�DI���mR�C���Cs>.E�|$B�=x�bAz�    I<�����1�Ţ�8E    %��    a*C���DŒF�;��C�F���N�o1���}�D�_��l&D��D�T���WFy�vD6�"E�@D�=C���Bm�H@�?��D}X[E̗�Ę�xEZs�D�aE֋�<�����Dk�E    �A(�    �4�EZt��(ID�<ļ(�@�(�wסD    j�D{D��&�_D��E5#QE&�D=�0B�y��}b*E    T�
�    ���C���B-��D    mF����ųuŰ��C�����jE�tBP�Ŏ0�E    �l�Ӧ�C    �&�CU���.�C���Zq@���p�K���u$E18C���CS��EI4B�K�A��D$S��5��D;�+�)"�w��ę����E�Cn��m��E,�ŠuF� ��Y��T"E��QD�ſ�Ĕ:Z�    ���B    Fg�WO'�L��DK�jm%E4�r��p'�Hx��yRBC��B��X��D|�J�?�.��e�-:D�c��A�/���'B/ξ���C�~�ſ���nlE    �>�C�Ų�Jg�    ���C±�D������BC�V��N-%ŁyB    7��C����(d*�C{eũ�/�!��<7D"f��,�4D                    *�aň��klD�����&D/�DQ��C
kD�k"Ħ ���D��\��c8��t0CAc�B�#n� �v��2EB�B�Ί����(pDD-Dwy����E������D�F��÷��q0DB[�Bl�-D��FG���'f��q:«�üY:C����^>ĂՊ���LE=+�Ì�)ě��E���R5�����Ǩ�s%Đ���AD3�6�D�ٍ�e(7E���C<s��2*��[��N�        e��z�%��P�Do�oE���e�LE���\����E�̴D&�m�ǢD���h)œ�OE�R�D�X��,G��x�wD�khEsS��CC	Z�C%CT,�    �AE׾C|�(E,�����K�m�c5(E���D���D��KDp�D�B��&��E��K���?Xę�E�=Č�B6�-D��Nđ��qx������(�E���=�����B�B��&�5��P^ĘF�C��J�*��D	��Cf�	Ŀ;��;��?��C���Dz��Ē���_���0/��2��ďd�D'���ER(D�7�ī������4� �l�E�aAT�EmR���GJ�    ��'Ņ���    ��E��<E��5�0x�š` �Jb{D�1=E��iD\�-�P�.Ļ�DU��C.�E$ ��!Æ�<D��ũ�pªPŶގE�m{BJ��ź�DeEd�D0�Bw�4E�������Dvg��G��D����'͋C��B�l�D�!~�    ^]E� �. 5�Æ�ž�U��cE#�1ņ�İ��:Ȭ�����D�����E|��D}E��DUpKĺ|BŬ�,E��E|��B����nè�4E�T2���E��}EE��y�����+��CpC�]qsD��l�    �g�׺DKhE�B�U���.��ࢉÉ�Ü���BN"ũ��}���(���P��D��0���D���D����)�D�.�DI/E��E    �"E��>E'p�D��Ʉ�D��.FT���G���u���
��Pr���#nC�C��D��V�    ��[D�DN��`DT^�E֍�D��Due��-��a��D"ȯ��$CB� ��7�BD0��C�$Ir�;'��1�8E��ĳ�BD����d�D^�Č���Һ�C��E/�C�5��͸FK^�r_%ŭ��D*LE �ı-�C�U�D��bø�E�pDC8�Dy�F�'�<EF�l�>��Y�2E�]�Է?E?y�C��B        �ݬDܨ���"�    ��kE]s���8�RyEv�!@��COM>D" lE���e}W���d�H�[ô�"D�1<Di�D    9�	�1�_�b��E������B!;�D��D�Ř�3��M����DGˉE��zD�D��DC�vDF�I�g�?D�#�Ee��C�I�IE
Q:�E!A��r��E�R���E���u��zDh
zC��o�p��Ò��D���    �rC���,��DYC$�K�E��E����:D        ���D�D4j�DJߍ�    �^��/�C5�C�Ҽ�P��DI]D�ۢ�2YBd�E�*D�@@E��������MD�� �@nq�`1�ė}�Ī5�D�)s�p�E�1�D�$D�!E#XD���'�L���E���D�ۇC��Dn��F'C����<{lCH,�� �ĵUFD�/E EQ<%<^E:5�D�l<� 2#��q|�/f��CQ�Ŵf*D�M�C        �E:�$C�S��
0)DG���$�ԦD���D����kD1B    �IGń��C��ÞJČF�D��"ŁA�C��`Di��B��%E��W��;�D�K���IBDTZ��    �;DV&�����.E������Ž=?�    �� �b���{ ;D���Ře%E�/�DrJEl�bE���B._�DFy=Fڠ�D    �V*��4r�bX+D���<Q(CTe�B�ŝ�,	��Xf�EC    A�^C�'E���E��	 �C E�#�D ��Cu?E<��Cz��D<�7�9!A�/���]̚�/��D �C_`IDӶ�B|Q�l��B����̑C��;E    ���D    �tHŀ�[��PdE��D=�#��A�D��C    E���U�7�lL�Ŀ�?o[F��Ņ(����;�8u��U�@D�=�Bx!��    n�9��@u�
ݏD&�ND����A�mEt���kz�D�sD��QDiR�3�D�L�DbM�D0��E��D���A_�N���{EbOC.4E'�?Ca�E�E��D�	�	E8	rDNȔD$�F�Xdż$,Ö�E�fE��D�t�b�n_iter_�N�
intercept_�h�scalar���hC���H���R��_sklearn_version��0.23.2�ub.