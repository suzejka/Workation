��       �sklearn.linear_model._ridge��Ridge���)��}�(�alpha�G?�      �fit_intercept���	normalize���copy_X���max_iter�N�tol�G?PbM����solver��auto��random_state�M��n_features_in_�M��coef_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KM���h�dtype����f4�����R�(K�<�NNNJ����J����K t�b�Bl  ��:3	M6���D���:�ĥ&E|���Q�����o����C�D�h������9�oň��ŦeFD%F�\*F�:�J�Ž-��,$�ŏ�A�K+aE    eX"E�Z��    GN4��NsF֝iD:���M�����6���M�8E6o��1�2E�h �t�F�b�E�9EC�I���}E������B�B�F�
?Cc�EE-�E�=�F�.(ű�T�    � ���"v��E����Ջ�Es�Fyn4D�&DC��R��8�El��    ���    '��E᭵B    MҘE3D���5��>ZI�:y]E��E"��DɁ���Ř=����Ds���*�E�k�Ñ���w��8
E�]��m�M� F�`ID�K��<�GE����f�D�~��Yb�D�[�Ć�%�K�zK�C�|;�Et�U�;���*��ּuD+�E�-Di�%��CT2�D�V�E�(�D�Jo�Fi�E�'�E�/R�.�� ����3�BME��SƻRrE�rC��C�x�Ņ�hF�;�EK��DN�E���E�\��svIƵ�+D���F��DǥE~Ѱ��Z"E$���    ?�ļ������D���T��D���E)�UƗ��DO%EW�ř+PE;�D_��K�p�GD �E��i�[�E�E        u�Q�2k�N�D    v���    �e�+��E    ����    H�7�¹�D���À��y��W�ļROE�ՉC�"��     �ËnDH$���fD�7F�A�DL�    n8��>��Ƈ���+tE;�����D�)�D��2D�H�Ġ;�DM"�D            H��D��D        ��@�            }��� �4E    e���׃����]��D�h������    ���    �b�D��    
{�Ŷ5-�    �ϟE        �v�@��ñ$���        �N�D        [� ė9XC���E    �v4�    o�p�        Y�C            �d��B�éDG&�ħ�m� K��    E�Ĕ��D������Et)}ō�zE�E�oUŁzM�B�Do��4�VD    ��y�L8DE��M��\�ĸn�ŝ"Z�=��F��Zœv��i;��%*�7���#�EQ&�i'C�´Cq�EE    %Q�D�ЀE    �0Y��lE�ZE �E���E���D埆Ù*/ŝ��F!��    �+�CoΖĝ �D��aET�����ET��D����yb��    (M	E    Ҥ�\W��m#�� �E��D    ���    �2b�<����EzLB����Ћ�����    �mJ�m�(D��$C    U)0E���iC؂lC2���L�eE    [PE��EX�X�    H�D�%F!bE��DD    [�ĩJ�DB�CC��D���            6�Ī	�D�<���PyB礪�    +X�D                �#<D_�=Ů�����E *T�    )ą�    U9�Cv�Ŝ�0E        ���    ��$D    �j~�U�Ę�f�s^D�<C�*t�L-	FmD�LEDr�    5�~��";����D����j5E�g\�s� Ex�=Ä���]��~�LD��
D�d��3�he�C��Û�"�\%�E���IŊc�����1l)�    زĪ��� E    G�4�s�C�����Q6š^�Eb��re�D0�t���SE�E�^�B��DHT@�    �<T�&��Ÿ]�        ?�E��4���C��Ē%����BY�]B�F�
�    	�:B2	DK�E    #5��E|�D:��D�U��    ���DK��r�2F��.�2��    �Ř�����?����PC�mD    �s�C�`$�S%�ĐC�D���DC�I���C\ٍ�    m֓D�zvDM�`ŉܙ�ח�����D��    C��    Z�>�)\XD    �L��xuQD��EBD�;�D�jE�ُ���D~�8�        �|[EO�D�K����        �E�SE    [��2���Cf��D���E    ��DTֆ�؆D        C�Fw=�C    ��Do�E��
E        �(E�E`�    C�DHdE        ��E    x��E�	E    ��-E        6{*�            ���Dc���    ���D��"�~h�    q��D���������]DL��y=;��.�    ���F�ÊA:Dc��E���DԨ%�    ؉��    ���DFY/�    ��D        ���ƥ�GE��[E��Ez�D��C���D    �`��f�\��D��a�N;d�d����y�A�EEDM��X�D���    a��        !/�    }���.R����F�G�D^�_D�6ƃbŜVE    1���j?;EiC�A>E�l��    �������!�E�����_�wu������l@B�|�������-�=�        �`D    ˋ*�L��.Ģ\�D݆�Eժ�ĩL��    ���BLv��v�ś>Ū-N�    Z��E
���E���{+FE    �E    *u��-u��    ���,��EJ�C�9��     �D`F��B~����EU2ī��            y��QS�D    ω�D    � �Ľ%B�$!aE        ���*oE�nE���}E�x���o��    F���D榡�D��C$N�Dx�D�-��G��D    E    ��E�4��4"D\9�E��=EZIŖ�kDAS�D�8J��0���|��[C;)��    }��E�_�D7 ���a�    ��j�ϭ�DoI�DtY�Ő��    0L�    �x�EoG����Ĭ��DOn�E�SE���EῨ�    Z��b��şFEk�YEbvfC�~�C]����DnW��@)WE�U�F0v��    H�E�KC����5J`E	�#E/�F1��3��\ZIE�,C    A[KE2�D    ձ�E�ƚ�� �C        wgD%~�C��A���    ��C6�3�9�7C��[2��dB            ��!D,��C����S��0��D]h�ɥtE�ecE        ��D9O�D�&�        ���Ĉ݁D5.�D    ��D    ̒M�-9w��.(�            �/ E�8 �|zGE�?�Ĺ˒Dd��ċt
E�%+E>�.E    �@�E���B����a���&�EJe6E    �U��`T�C�K��1��    0&�5��    �1��ɖ�E�[��q�r�+OD�+�tE�ŝ�!��A��<߃E���C    m�C��C    ��C)���b��E�k��    `�>E    ��SŰ��E���    �M��ODmE�.�D    ��C''�F    -��|�Ƽ�UE���ăE#W+E#NFn9"D�Jj�W��EQ{E��D���ʂ�� Ea�%Œ�3��4��#.VDe�@gw�    �E    �����-E�#Ei��d��E�SjņN���|�$�jD�{D    ��:EX��    �=D�����k��    =�Zū�8D    ����96���D����    x�F�>E3W=EG���    �N��R>E?��E��MCL�aE=��E    �hD�b��    V��|{�FI��E��~E�����]~D}�Rď����Bn�AT&�    ���BT�1�        �Ű���            <����p��D�V�D#8�1�l��rC��E                V"��DIů� Ep���V�EZArDkKE�[�D    ��*�'�����D    6���]sć��D�&eD��j��D�P!Ea�� j
E~��    �bZD����    m��    O4X��	F��%E    "�<E    ���DMn�        Iޏ��{E    %�CC    C�D����    ��E�/��57�V�/ņD��    �"��        �&��;5J���CF��z��Z�D3J �m}���     ��    w N�    �=}ES7F�r��E    ��F�K����E��    }��    ������FZ��E8\�Eo��r- �m��E�<��4�E�	�ǘj�9�ŀ�SD<�F{�G����QN�4z���Z���|F��DZ*��    ՚a�    !AF��DÍSE������    	>��$�+E�TD�[C�IaÛÁ� �E��*�     JD�_EEJJwEH��J�C�Cĳs�DO�aD���D����*��^�&p�    ��rD���~;��00�C��Ø� �x��C�@/DID�4B̆���ŗ&3�<�E�4��˜�D�DESL�    �����E�\�R��B_� E~�D#���>E����=�D�݋��Dn̲C"�E�fE/]�E��#EML�DP��C(�E�<n��tE�ICM�DQ�&���c�naE                m��E�.G¿�`�cS��I�E    ��ƵفD�%!��s E&eC��    i�K�    ���K֐��2D'�
�s�C    �O�    e���F`��.Z9E��E���Dt�DnJ	��D�ڨ�D�,��0�]�6D��DūL�W��D�EM/D^E�C�%
EB�C���×���L/F8v���XŊ�D;.�Et_/�!!D4��;0��YrD[���ul�D�DB�V�D�=E    �i F��D    ��E�3�C���á����0gĝ�ZF�C�4���J��}m��g��W!E5��D��ņ�i�"�E    �1�ğ?�D�YE�/�    *9�Da��B��D<J�    ���D�MD�,��SE�Ss�n�����T�=@�dQ�CJ KE    �GuD    ����{6�D    �a�C"�.�O/L@���C����EC&ID�D��yE    �-AE5ƏE    b��D�o��0	�C}HfD,��E`�%�F`����s_İz��׾�D��YD�EO�
E�DU�HE,���[CE ��ĺ���U�@�ب���"tC�7��"Y�r���6%3�0��ĳ|/E|�D
w�Dz���    ��'E    ^�-Ś�&����>��Ŷ��8&���A�uIĨ�ZEz��D��b��dn��+ĮgnE����f(ņ���y�C}�ĒI����;�/D�,�'z�E�.A�ߌ��H%�C���D@C�íz0��?�����`�B����g���U�D    5�E���X1ŭE���ĎJ�    ���C    3�jì�!D,@��dō��D���C�-�D�}��շo��F��N�D5R4D�]�D����>D%|Š*�E�d��d~�����M��Ȭ�Sň�DY�\��G��ϓ�Cr�ů˸Dؖ�DB��D̅D.���s�JE��E�.�D����{�D<��&veC��pDE�5�C�ͮ���@C+��C\�����QE�e�Ç}E; D2��Æ�AE���DA�����D�JE|@�4<}Ċ:E�^��WE���qDk�]Ef���M�B�fV�B�r�E�%@�։�U�E��{�6��C���C�%V�4A�DLCMEM
�#�C�����R8E>^�D~v������1��}�EE�D)fd���K�    ��uE�N����-ŗ-����@K�Df� �U�į��C��E    ��b�F5(Cl��i���������U��Dj�C�:����б���E�D5�C��D�uv���D��C|�3E��Dn���3C��D�HfD���^�D� CEμ%�_��Dv��8�x��[rķ��÷SV�[��F�:�&�ǞDT�D    ��<�    u�5�1���|�+�$���Ɯ�Ġf�D���*Q�D~OD����!EC=-�2t��/����yE��C��&EA#�Cs4\ĳhN�q�D�8�É<Dpj�ą�_ĭ����y��ĊI�:���V�Ń�����EO�Ē.�D����A��)E�1���p��gD�k.D2[Gč�G�2�D�LŹ����D��IE36ĩZA
?�DR��D�E闃�˘��1>\C�h��%N�G��ӮQ�:3��ģ�p�[���/�uC�	�ģ���G�D}�)ňS�Ey��ĆA��Hn@D�k����DY$�C7��Q[�;"Ī���[�s���$DZ�/ķRG��e�C�t���Eħ�\DЁ�D�#EσXDZ����1$�R�DYxDv��`VsŪ�1BMoj�!�$E    5vDF̿�;�Da�7�Y.&�K`���D�$ EF���ĜD���v�ê���\�k��ǯ���SF    BO�C¯a��ˏDipE�QДE�S�Dt��_	����cE���W�B����t�����DF�SE�MQEt�EkDe߇�Q��F�i�RE���/d1�`�2D�F�'�E�OE�܂ĳ�_D�9�EXuCD[0�ð�(�7��C��Į�Y�I{E��J�@�I�^WMD<D���M8A�    ��;C		YD����D�Z����Ş��$�E�����5D��0��b�C9�œ{�D�B�E�nF��Cr(�h�?�8)"D�kSD���ĝK|Ĵ���j=�D�vD�`�B;׎� N
�v�Ŧ��DS�,Eh&]EM��C����C@�<>p�dj� ��s��E&ѫó��D/T�ġ��D�� Dُ��o3wE?r_D�0�Dv��/7�B��!�LCE��E��LĆM-��	`E    ��D��VD5F�.�oEw��EtLFES���:�%C        ��ŋI�DFV�Cs	ń���cRD    d@C�|��fU��I1���q�D_���Ɔ�B�^D)*�E� RCE��DB��D;�mDVW�i�4EL�B�    �W���E�t�D1��D�%!��e�D�P*����Ĥl��    �1HE�2H�    �E��7�;Ł�CF��DDC[�Co2E�:���'��lpD��.�y^�D>�$�ec�C�0�D�����!	MD        �����*Df�x^KļD���;��1L�ĭ���&��    �E^R�CPH�C�����C���JƽD�uc�Vc�P���_��C}LiÀ������oEq� ū��͞�C+C�D�����E}���	ìſD*�Ŀq�DsE�D����i�-E�	dD`V��+~���s�EQ�?C���C��BW���**������U�o ���D��U�    ����9�C�g~��5�E�7���A&�U����I[D�XD���Ĥi���RiC5Z"C�����D��+��6�y��D�fy�z�]E�Fś��jB�s]D�eL�                    S���Ō6Ep�`ŞE;�Ϧ�D�#p�    ��wD        ��������D�D    ���D�XE9�7E6�S�A�kaĪ�nC    ӋaD�ֻľ��D�hD�ƵD�:C    �UxD�4��~"��Ȁfč41ĶtyE}��D��En�Ā���"�0�b.�E��B�ęä�8E���jјDZ)Cſ���n�$��2��`����DV����NnD�
�İ"�B߈"�O +�m�^š�xĔt�b�n_iter_�N�
intercept_�h�scalar���hC��I���R��_sklearn_version��0.23.2�ub.