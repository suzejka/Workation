��0       �sklearn.linear_model._ridge��Ridge���)��}�(�alpha�G?�      �fit_intercept���	normalize���copy_X���max_iter�N�tol�G?PbM����solver��auto��random_state�M��n_features_in_�M��coef_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KM���h�dtype����f4�����R�(K�<�NNNJ����J����K t�b�B�  �O<CĻ6&'��z�ă�6DzaET"��Tk��&�Ĉ��Du�D�k'��x���SE�`�E\��$�'F�E/��:B��E�/�ĳ�����E6tOE    �G>E�'E�e�E�ũ��En�D^K����C?@��E���sYŉ�L�    ��pE�QE����$��CK}Ğf�Ł��Ã�E�L�E���ơ6��kE    *�D�cE�=�j4�E    w��D�I��o��D�ȏ��DE    eq�Ż�>��6"E,��ò�EEJ�E��D��e�3e5Ź|�ı����8��C���|����FŲ	Ũk�E���š|?D8E�ŀ��Ei���|uUEj��Eo����C���EcyUE�N-F�7E�c�E��TE�@�D��ƨj�-�    ��pE��E4� EG-��Y�D	�E��D��'E    ,��-�Ea��D)�o�D�h�?F�e��.-�S�~E-�ZDi~�į�^E*Y�BcL�E$���OF�b�EǋTEǍ�Ab#��v�F��E�>MEï�Ƴ;�DC��ũ
2E3_��8DE���D    f��D��ź��ŉe�E�������HV�D6#-F5�QE    [�d�    \
AE}�������ň�Q�;C�C V$��*)DT�|E�^�        ��A���À�D\E1�
E    �x>E�%�E�m������        P��D�Z�ľ�Ĵ�iŲ���3y&����prD    ��@D� Ŧ˩DxX���:F�2D    #S�`äE���FɈŒE�J;B΍D����/�
D�<�D�4EV��        �j�D.��C        a�C        �XRD���z*�    P��C7�Wſ�Ħ�,EƓ�E    w'�� ��ĝg��"2�Ī,�A~��]�5E    ����Rf��    3E5םD���A����    :��	�cD        k4H�    �/�    ڞ&E    ���D    ��TE���DO�D        wLŗ�J�    {*A>�EjRC�q�Ť�&�ܚ�v��D�@�������CV�;A�C    ��E�;�    E'D[��D��qũ<�{�mF�R�C^����#��?���E�D&�_҉EНE�Y��    �κC�D��,�k����C.j��&[qE        �
�E>M�6ζ�)��V��;HE(��M!�ߋ��    ��D�;xD�\XD=��    B�D�b���[�����z���lE    Q�#E0����`ŭ^E���D    ��Db��h�'Ep2>Œ��DK^D�?BE�G>�^�D    yv�D�����/A�    )�Ĳ!E�p��E8�B۬�ŔT��        �ǫ��]
E    C��C�I�EK�dE���C    ����O	�ĸ�B	d;����            ���BY�D�����Dݑ�D/�`DP��ĺP�D            Ϻ�Ck�����C�E����    ߙ�����    ��FEW ś��    ��%D    ?3RB    ���C    /�W��\C�[Y�$�́�
�vĐW�
D    �xF`M�C1�����ŉ(EZ��U,�D�J ����9q�$���/��B�Dv9��J�.D�:�Cm�C'�ũ|bD.�8�| ��2�'�����    ��D���Do �        &��B�ņMAŁ~]Ū^=C�D�K�  O�    ��LC��EԻ.E    �C�.�E�-�        ��4E�7(E-FT�Ņ�9D    ~r�ѡ�E�g�    ¶�B�!C���D        �oD�j�đۅD    |	�F��Ė���_��D    �����PE�ۈC���Ž;aD��D���        �4���D    �y�CCTŞr�6��DX�x�DĻ�D�ޑEe
E�<�N��Bp�ŭ���    G��D�AŖn.Dw���֐D·�EޮE�c�D��3E9�D?>D�$�E        _`��52;D3=E�P��        Ì�FݧE    b�|E����hD    �	��$[)��p���}�C        �|�F%52E    ��Dd��D            �!Ź7�D�)KĽ���        ���DtK�E    �X�����D    ����t�YD[�K�,�D        O�	D_=D��    W���W�]E�JQE    %D!?�]-���Ŵ^���ݧ�F�*E    ���D/S�J�RË��    ��h���    :\�Ę�(E[�4�g��D        p!�ŘoĐ%h�ĥE瑶D$r0��b�    ԣeE���ţ)�ߦZE
�yDgV����+C]��C��E��Ŷ�b	/��d��        ����0�D,u7��P��I�[x�a�EF����s��C��E    '
�Bs�D    ���DOu�D    ����á�D!�\E���b4H��`���EЌ�D��aE!���E        ��C    ��KD�|Fc9��!U$Ev�ŊVD����	�@�    ;��U��o�>E�O�D��D�    �Ylİ8@�    ����_F�8 =�    ����    ��D�|����ò8��    ��D�J(�"
wE\U�'��D    ��aEݘyE�)�D        9*�A�%D    4�oD@�������0E��RŎ�+�        �;7E�ؐ�+D���    4z��Z�s���9�Į�c�{������E�iAEo��(�N�
��    ��D    f8�ĵ!s��(x�ťVElq�Z�E�� �˔�D�@_ơ2�D    C^Cr�E    )ֆESk�D5W�CM��    ��/E}�Q�%�gD�&k��"D    2��    vbƣ�E*�Zň�i���2����.@=�^��HI"D~�D��U���E��Db�b��DɻJ�P?�U�DԪ�S�>EZڶF]"��    #r��b�wč~J�(7�D�    �%�D�'�g�:�eE�C    ����C�o�E'_�E,N�ܴ�D�i��%�-Ñ	��)(�ķj�
�E    ���Dň2E�I��R���~t��Z�C            �uY�c�_�:$#��p?E��D FD'Bv�
a��        ��)�.ܼD&�A        "�7��ƌD���D    ���*U��	���B�m��yE            ���D    �"�ĉi�#GlD�?��    �B;�ZE    �|�;��Ĕr3F�����ƞbN� ��Et���n�DD� � ��E    ��!ŏW�Ŗp�C�
fE+���*�6Y���w!�	�^�S��D    �i�����Eȴ:�    �/Eqa�D    V�Cׇ7D�l�E        ���4��C�я�{x"E��D    �l���[�E��h�)׾��z�B~2 �    ����jmF��;Eu�/�C� E�-Ec"�E&����,�e��J�^Ez��A�B��&͂D�E�-�}�c�    ��D� �E-0]FЇ�BB�E�    ȉ�    �Z�x�E��^Ž|2�E)�E��=��
EWl��    .��#>Eo�/D    �&��7�]�于D    ��ME=B� DįSDP;?���R����zű9WE�HE�X9��AfE    �Qť<E\�f���
D^\?śozE    ��a�x�>�    �kE    0	ƶY��.@9Ec��&)C4�8D    �E    X�ĺ�0E        ��fE[��C            E-Ĭq�C��V�_��Rx��,E�� �G;��                ,��ŏ��Dl;�Ċ�}�&q�E[��ď�E��D���E�����2�D    ���Ds���U�FD��D��OE�����z����A�Dd��D    &s�C�UQ�    2�$E    ��nF&(Fv��D    �x����E1�D`��D        A PC9�EE    ,!�D�'�D�����s�E    ~�F��]�ȍ'E    0��Ç��D��QE        b���F+E.���K��d�@�h����B�D    R��I�E    r�IG    �l�xv�F�F    $��ł�=E�|`E�!�C    �oD        ���F6��E YCF@^��qI�œ7��a���vO�õr�rC��Q5*�X�yŞ����y G���ÙpWE���d��E��6��N�i�m0LŖG�C    �}M�m�;C�]���5�Ś=�� ;D�    r����-�a����wD��7D��E�R���U8�XC�ĥZ�ÔN?�����U�Dŷu����D�ĳYELwE'���4E�.2D�slE��&�*m�CT�"CE��C�^C� D�e�¤G\ĥ�n�.��D�+�����2�k�m��Iў�hoyD"�DD    ��"D;��^jc�u;��%cE��E��D��D�)}C�Ċ�BEt?�E
����pEXo\Dw������G��D.U5��A�E�d�P�qE>�-C�_���IEKz��n;]CUl�D3��Dl8(D��
D31��                g��E�F���C42���$�D    ��#�}I�DE����/BZÓ:�    ��,�    �&���qC�p��Bx�y���    ��R�    �+Dr���    �1��܌�C&*�D-h�C(��D�XjDp����Dċ�C!��E��Dt�E��Emܚ���D��COt����E��)Dd�o�M��E�lŇ^_�    `UxC�aeE)���� ~�XF�ĵհ�P���G�D�a�Ă�EI�WEvF�a��    ��ō�Y��x�{sD�mCBQTF�0��YD�ĺYME9��B	���@�D�9�D��D�*�Ow5E    ���CM��Db�IE��D����!T�DҼ Î��D�4��      �C�6���:D�FYŞ������ŁePD�DCL��    ivSE    �Dd�D�X�C    BvQD�=�D�Y�CŨX�dE�^��h��i���=*�E    W�"E���E    �EG�fC}\XE�ĸ�\E|���E�n�DCh�{
C)o�Ī+��-��:�`�D�*�Ċ�D��$E[y�������Q�ÿ	�ü�����E���m%Dgr�D-ׄDC����Z�D        �X��    �SE�)E՜�Ė~�Ō�DE�B�UC��,�+�~D-�����˯�;1�+*��	u E;�C�<���V���/E� �C����G/ĩ ���6�E    ��i������ñ	��4,YC⍅�o�Cs����E70�    \UD�W��K��CD[��]�g�g�����    ��v�~"�    ̦:� �Ħ��C    �@JŠN�D�K�D	�]��t2Ĕ�D�L�À�.�2�C:��DwT�D܎ C��D8�����r��Ŋ]�Ê��B�[/C�/DXX������DE~OEIhJĽ����%E)+Eu(��J`ŮV�D�W�Î;F>�D}���vf�D�˞C��5���]X�    ��Ch�uE]���kʫD�x��T��D����J�DGnbEEH"D��DT�-ŖA(�� hBy�2œϽ���D�p1Ŝ2Ɣ��x¹C��!�ၑC֚�BR�Djw�Ÿ��Ď���y��D�ZE�R����j���-<E�Wh�(a�D!D&�og³�j�RD�R�ĝODě1)Ÿ�xD��ADӍ�B4T.D�0GE[�m���1E�ƃç�ŉׯD���DS�l�.j�����ÃȻBŷ+�h�D��D2=�h��Ċ�hD�҆CU�d�B4�C���CEa�NēU�DZ���S�o��6�E^�C�MDL�
Ă@�D�VaEҔ�D��������}D�����|��uND�1C�RػD�-��t��DE��㚪�8t+E�G�Ē1U��
�p �H��k�    g�ġ���    ە�D�_�Db �Ðdń&D��D{�B�8A$������D�&�E��D�XJE ������?�Ŋm��!��D�mE2����D�#�D��$��שC�<�Bm!QEJDcD�v_C���!��z	�3��EH�Đz�ōڕ��EE5��ݓE>�&E	�;�W���r�k�^�ě��D|� E        �S{�a�Z�    3��C��E����+�D�E��G�e{��y�D�8�� �Ég�Dp��C�)���KEiw!��w�Ú�EE�{�H�4EgkC�RWï[����Dp^C#J�DX��ā�D��%�5DN�Dq��DţI�ڑ	ES#��g�Ei�>EP~��ˑ(���D��C�ۢC��ďb-�6�D���� �E��$E����۵OŘ����ĥY&EŃ
Eg���҈�D        ��D�yDfP�N�E�*�e��DUX�]���	��MʮC%.��ɂ����uF    ���D?ߟ�֢�CJtE��o���ħ����Ġ?�D�ЧĈ��C�ùD���/H�DB�( EAԤC�`6Aބ��o���    �{��� �Dy|����DNW��Un8E8�����gE �8E���$��B    &ӄ�#�R��D����<���E�����EE٥"���2�݈�¼��A�[E��Ũ`TE҉�?��X�9�    e��`��C|�Ń@�F    vu��N~Ewv�E��D�BE���(��įL���ljE?��[D7D���ó�~Ī�D�4��)����rE����%N~Ü��    S��D�7E����j��nw��h��C"�D�H�1�tD��Do�����ME�����M�l��DKh��Ft���$�D�h�š� ��d�D�i�Dg';E�K�CI�+C2�^�C�Tăh6�    <4DY	E#1�D�bE��4E͋&ń��Dd�D        ���В�z<UDK�D��A"4NDy_��}�RCM��5P��{�D��CI4DC�y�o���    ��D��C%:�Df߁E�w+D(�yDh��ŠEҥ^��}>�.MD	3LDtE���Dv2E� �    b�9E/\xD�� 4��c�ΠpC�oE��B�F�D�pC�v7D_����B�E��]�ÿ�C"A�        �"��/����Dd��z
���D�����9E���    �7E�þC����rf�Ø��ğ� ��gD�>��I��C���ğ+���C~�ů�7D���D)��C!��D ���    �	D;��Drs��#ϑ�-"�E,x�C�/�D[wĆ�[D ��D���K�D)�A��E�`��EQ��0gy���D]�D�'�Ħ�aC��3��cD%^E���    J^�C3��C    e�C���D���ô(�ŉ~�Üp�ó�#�̉D\aD!,D�:�D24��.rPë�Ħ�pD���D�B D\DW�(E�����[D䐎C��1C�o�D��(�*��B    �\��    �kWE%��A�R�T)����D���D���        ��C��@1_��M��8D��$EXZE����e������A^��    �e*C�pC�$��T^�D�,�    ����a=�$�D�h�ľ%D�	�D�i�D�YŤ����o�C݅�E�!�CI��D    ԄE��#D4��ۣ�~ EEq�3�şܣ�*ڦ���D�ǥD��6EsD��$D�<IEmP�Ĕt�b�n_iter_�N�
intercept_�h�scalar���hC7�
I���R��_sklearn_version��0.23.2�ub.